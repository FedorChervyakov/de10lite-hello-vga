library ieee;
use ieee.std_logic_1164.all;

entity hello_vga is
end entity;

architecture A of hello_vga is
begin

end architecture A;
